module RISE_EDGE_PULSE_LENGTH_CONVERTER
#(
	parameter DEEP_PULSE_LENGTH_BITS=3
)
(
	input 										IN_CLOCK,
	input [DEEP_PULSE_LENGTH_BITS-1:0] 	IN_LENGTH_OUTPUT_PULSE_CLKS,
	input										 	IN_PULSE,
	output 										OUT_CONVERTED_PULSE
);

wire OUT_SHORT_PULSE;
Pulse_shortening_device PSD
(IN_CLOCK,IN_PULSE,OUT_SHORT_PULSE);

reg	[DEEP_PULSE_LENGTH_BITS-1:0]	REG_CLKS_COUNTER;
reg	[DEEP_PULSE_LENGTH_BITS-1:0]	REG_LENGTH_OUTPUT_PULSE_CLKS;
reg 											REG_FSM_STATE;
reg											REG_OUT_CONVERTED_PULSE;
localparam STATE_WAIT=1'b0;
localparam STATE_PULSE_ACTIVE=1'b1;
assign OUT_CONVERTED_PULSE=(REG_OUT_CONVERTED_PULSE|OUT_SHORT_PULSE)&(|IN_LENGTH_OUTPUT_PULSE_CLKS);
initial begin
	REG_CLKS_COUNTER=0;
	REG_LENGTH_OUTPUT_PULSE_CLKS=0;
	REG_OUT_CONVERTED_PULSE=0;
	REG_FSM_STATE=STATE_WAIT;
end

always @( posedge IN_CLOCK)
begin
	case (REG_FSM_STATE)
		STATE_WAIT:
		begin
			if(IN_PULSE)
			begin
				REG_OUT_CONVERTED_PULSE<=0;
				REG_CLKS_COUNTER<=0;
				if(IN_LENGTH_OUTPUT_PULSE_CLKS!=0)
				begin
					REG_LENGTH_OUTPUT_PULSE_CLKS=IN_LENGTH_OUTPUT_PULSE_CLKS;
					REG_CLKS_COUNTER<=1;
					REG_OUT_CONVERTED_PULSE<=1;
					REG_FSM_STATE<=STATE_PULSE_ACTIVE;
				end
			end
		end
		STATE_PULSE_ACTIVE:
		begin
			if(REG_LENGTH_OUTPUT_PULSE_CLKS>REG_CLKS_COUNTER)
				REG_CLKS_COUNTER<=REG_CLKS_COUNTER+1;
			else
			begin
				REG_OUT_CONVERTED_PULSE<=0;
				if(!IN_PULSE)
				begin
					REG_CLKS_COUNTER<=0;
					REG_FSM_STATE<=STATE_WAIT;
				end
			end
		end
	endcase
end

endmodule
